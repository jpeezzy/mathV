//GENERATING  A MAXIMAL CODE SEQUENCE.
//MUST HAVE 2^n/2 ones and 2^n/2-1 zeros
module maximal_sequence #(parameter CHIRP_WIDTH = 1024) (
	input [CHIRP_WIDTH-1:0] in,
	output [CHIRP_WIDTH-1:0] out
);
	always @* begin
		
	end
endmodule
