module fast_inverse_sqrt(
	input real x,
	output real y
);

always @(*)
begin
//Begin the inverse square root
real x2, y;

end

endmodule
